module tb;

// IO
reg		clk;
reg     rst_n;

/////////////////////////////////////////////////////////
// TEST
/////////////////////////////////////////////////////////
initial begin
repeat (10) @ (posedge clk);


repeat (5) @(posedge clk);
$display("Test completed");
$finish;
end

/////////////////////////////////////////////////////////
// DUT
/////////////////////////////////////////////////////////


/////////////////////////////////////////////////////////
// INIT
/////////////////////////////////////////////////////////

initial begin
clk = 0;
rst_n = 1;
end

/////////////////////////////////////////////////////////
// RST_N
/////////////////////////////////////////////////////////

initial begin
repeat (1) @ (posedge clk);
rst_n=0;
repeat (1) @ (posedge clk);
rst_n=1;
end

/////////////////////////////////////////////////////////
// WAVES
/////////////////////////////////////////////////////////

initial begin
$dumpfile("tb.vcd");
$dumpvars(0, tb);
end

/////////////////////////////////////////////////////////
// clk
/////////////////////////////////////////////////////////

always #5 clk = ~clk;

endmodule